`include "uvm_macros.svh"
`include "LFSR_if.sv"
`include "LFSR_seq_item.sv"
`include "LFSR_sequencer.sv"
`include "LFSR_sequence.sv"
`include "LFSR_seq_lib.sv"
`include "LFSR_monitor.sv"
`include "LFSR_driver.sv"
`include "LFSR_scoreboard.sv" 
`include "LFSR_agent.sv"
`include "LFSR_env.sv"
`include "LFSR_test.sv"